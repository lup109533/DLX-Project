library ieee;
use ieee.std_logic_1164.all;
use work.DLX_globals.all;
use work.utils.log2;

entity FETCH is
end entity;

architecture structural of FETCH is

begin

end architecture;