library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.DLX_globals.all;

entity CU is
	port (
		CLK					: in	std_logic;
		RST					: in	std_logic;
		ENB					: in	std_logic;
		INSTR				: in	DLX_instruction_t;
		-- Special signals for TRAP instruction
		ISR_EN				: in	std_logic;
		-- Control signals here.
		RF_RD1_ADDR			: out	reg_addr_t;
		RF_RD2_ADDR			: out	reg_addr_t;
		RF_WR_ADDR			: out	reg_addr_t;
		RF_RD1				: out	std_logic;
		RF_RD2				: out	std_logic;
		RF_WR				: out	std_logic;
		RF_CALL				: out	std_logic;
		RF_RETN				: out	std_logic;
		IMM_ARG				: out	immediate_t;
		IMM_SEL				: out	std_logic;
		PC_OFFSET			: out	pc_offset_t;
		PC_OFFSET_SEL		: out	std_logic;
		OPCODE				: out	opcode_t;
		SIGNED_EXT			: out	std_logic;
		MEM_RD_SEL			: out	std_logic;
		MEM_WR_SEL			: out	std_logic;
		MEM_EN				: out	std_logic;
		MEMORY_OP_SEL		: out	std_logic;
		MEM_SIGNED_EXT		: out	std_logic;
		MEM_HALFWORD		: out	std_logic;
		MEM_BYTE			: out	std_logic;
		X2D_FORWARD_S1_EN	: out	std_logic;
		M2D_FORWARD_S1_EN	: out	std_logic;
		W2D_FORWARD_S1_EN	: out	std_logic;
		X2D_FORWARD_S2_EN	: out	std_logic;
		M2D_FORWARD_S2_EN	: out	std_logic;
		W2D_FORWARD_S2_EN	: out	std_logic;
		STALL				: out	std_logic
	);
end entity;

architecture behavioural of CU is
	
	type stages_t is (
					DEC,	-- DECODE
					EXE,	-- EXCUTE
					MEM,	-- MEMORY
					WRB		-- WRITE BACK
				);
				
	signal opcode_s				: opcode_t;
	signal source1_addr_s		: reg_addr_t;
	signal source2_addr_s		: reg_addr_t;
	signal dest_addr_s			: reg_addr_t;
	signal func_s				: func_t;
	signal fpu_func_s			: fp_func_t;
	signal immediate_s			: immediate_t;
	signal pc_offset_s			: pc_offset_t;
	signal op_type				: DLX_instr_type_t;
	
	type hazard_pipe_op_type_t  is array (DEC to WRB) of op_type;
	type hazard_pipe_reg_addr_t is array (DEC to WRB) of reg_addr_t;
	
	signal hazard_pipe_t		: hazard_pipe_op_type_t;
	signal hazard_pipe_s1		: hazard_pipe_reg_addr_t;
	signal hazard_pipe_s2		: hazard_pipe_reg_addr_t;
	signal hazard_pipe_d		: hazard_pipe_reg_addr_t;
	
	signal target_has_s1		: std_logic;
	signal target_has_s2		: std_logic;
	signal exe_source_has_d		: std_logic;
	signal mem_source_has_d		: std_logic;
	signal wrb_source_has_d		: std_logic;
	signal exe_can_forward_s1	: std_logic;
	signal mem_can_forward_s1	: std_logic;
	signal wrb_can_forward_s1	: std_logic;
	signal exe_can_forward_s2	: std_logic;
	signal wrb_can_forward_s2	: std_logic;
	signal mem_can_forward_s2	: std_logic;
	signal exe_source_is_load	: std_logic;
	signal stall_s				: std_logic;

begin
	
	-- INSTRUCTION UNPACKING
	opcode_s		<= INSTR(OPCODE_RANGE);
	source1_addr_s	<= INSTR(REG_SOURCE1_RANGE);
	source2_addr_s	<= INSTR(REG_SOURCE2_RANGE);
	dest_addr_s		<= INSTR(REG_DEST_RANGE);
	func_s			<= INSTR(ALU_FUNC_RANGE);
	fpu_func_s		<= INSTR(FPU_FUNC_RANGE);
	immediate_s		<= INSTR(IMMEDIATE_ARG_RANGE);
	pc_offset_s		<= INSTR(PC_OFFSET_RANGE);
	
	-- CONTROL SIGNAL GENERATION
	RF_RD1_ADDR		<= source1_addr_s;
	RF_RD2_ADDR		<= source2_addr_s;
	RF_WR_ADDR		<= dest_addr_s;
	RF_RD1			<= '1' when (op_type = R_TYPE) else '0';
	RF_RD2			<= '1' when (op_type = R_TYPE) else '0';
	RF_WR			<= '1' when (op_type = R_TYPE) else '0';
	RF_CALL			<= '1' when (opcode_s = TRAP)  else '0';
	RF_RETN			<= '1' when (opcode_s = RFE)   else '0';
	ISR_EN			<= '1' when (opcode_s = TRAP)  else '0';
	IMM_ARG			<= immediate_s;
	IMM_SEL			<= '1' when (op_type = I_TYPE or opcode_s = LHI) else '0';
	PC_OFFSET		<= '1' when (op_type = J_TYPE) else '0';
	PC_OFFSET_SEL	<= pc_offset_s;
	OPCODE			<= opcode_s;
	SIGNED_EXT		<= '0' when	((op_type = I_TYPE   and signed_immediate = '1') or
							     (opcode_s = ALU_I   and signed_alu_op = '1')    or
							     (opcode_s = FPU_I   and signed_fpu_op = '1'))   else '1';
	MEM_RD_SEL		<= '1' when (op_type = L_TYPE) else '0';
	MEM_WR_SEL		<= '1' when (op_type = S_TYPE) else '0';
	MEM_EN			<= '1' when (op_type = L_TYPE  or
					             op_type = S_TYPE) else '0';
	MEMORY_OP_SEL	<= '1' when (op_type = L_TYPE  or
					             op_type = S_TYPE) else '0';
	MEM_SIGNED_EXT	<= '1' when (opcode_s = LBU  or
					             opcode_s = LHU) else '0';
	MEM_HALFWORD	<= '1' when (opcode_s = LH  or
					             opcode_s = LHU or
								 opcode_s = SH) else '0';
	MEM_BYTE		<= '1' when (opcode_s = LB  or
					             opcode_s = LBU or
								 opcode_s = SB) else '0';
								
	
	signed_immediate	<= '0' when (OPCODE = ADDUI or
						             OPCODE = SUBUI or
									 OPCODE = SLTUI or
									 OPCODE = SGTUI or
									 OPCODE = SLEUI or
									 OPCODE = SGEUI) else '1';
									 
	signed_alu_op		<= '0' when (func_s = ADDU or
						             func_s = SUBU or
									 func_s = SLTU or
									 func_s = SGTU or
									 func_s = SLEU or
									 func_s = SGEU) else '1';
									 
	signed_fpu_op		<= '0' when (fpu_func_s = MULU or fpu_func_s = DIVU) else '1';
	
	-- ALU OPCODE GENERATOR
	alu_opcode_manager: process (opcode_s, func_s) is
	begin
		if (opcode_s = ALU_I) then
			case (func_s) is
				when SHLL =>
					alu_opcode_s <= SHIFT_LL;
					
				when SHRL =>
					alu_opcode_s <= SHIFT_RL;
					
				when SHRA =>
					alu_opcode_s <= SHIFT_RA;
				
				when ADD | ADDU =>
					alu_opcode_s <= IADD;
					
				when SUB | SUBU =>
					alu_opcode_s <= ISUB;
					
				when LAND =>
					alu_opcode_s <= LOGIC_AND;
					
				when LOR =>
					alu_opcode_s <= LOGIC_OR;
					
				when LXOR =>
					alu_opcode_s <= LOGIC_AND;
					
				when SEQ =>
					alu_opcode_s <= COMPARE_EQ;
					
				when SNE =>
					alu_opcode_s <= COMPARE_NE;
				
				when SLT | SLTU =>
					alu_opcode_s <= COMPARE_LT;
					
				when SGT | SGTU =>
					alu_opcode_s <= COMPARE_GT;
					
				when SLE | SLEU =>
					alu_opcode_s <= COMPARE_LE;
					
				when SGE | SGEU =>
					alu_opcode_s <= COMPARE_GE;
					
				when others =>
					alu_opcode_s <= MOV;
			end case;
		else
			case (opcode_s) is
				when SLLI | SRLI | SRAI =>
					alu_opcode_s <= SHIFT;
			
				when ADDI | ADDUI | BEQZ | BNEZ | J | JR | JALR =>
					alu_opcode_s <= ADD;
					
				when SUBI | SUBUI =>
					alu_opcode_s <= SUB;
					
				when ANDI =>
					alu_opcode_s <= LOGIC_AND;
					
				when ORI =>
					alu_opcode_s <= LOGIC_OR;
					
				when XORI =>
					alu_opcode_s <= LOGIC_AND;
					
				when SEQI =>
					alu_opcode_s <= COMPARE_EQ;
					
				when SNEI =>
					alu_opcode_s <= COMPARE_NE;
				
				when SLTI | SLTUI =>
					alu_opcode_s <= COMPARE_LT;
					
				when SGTI | SGTUI =>
					alu_opcode_s <= COMPARE_GT;
					
				when SLEI | SLEUI =>
					alu_opcode_s <= COMPARE_LE;
					
				when SGEI | SGEUI =>
					alu_opcode_s <= COMPARE_GE;
					
				when others =>
					alu_opcode_s <= MOV;
			end case;
		end if;
	end process;
	ALU_OPCODE <= alu_opcode_s;
	
	-- FPU OPCODE GENERATOR
	fpu_opcode_manager: process (fpu_func_s) is
	begin
		case (fpu_func_s) is
			when ADDF =>
				fpu_opcode_s <= FP_ADD;
				
			when SUBF =>
				fpu_opcode_s <= FP_SUB;
		
			when MUL | MULU =>
				fpu_opcode_s <= INT_MULTIPLY;
				
			when MULF =>
				fpu_opcode_s <= FP_MULTIPLY;
			
			when CVTF2I =>
				fpu_opcode_s <= F2I_CONVERT;
				
			when CVTI2F =>
				fpu_opcode_s <= I2F_CONVERT;
			
			when others =>
				fpu_opcode_s <= F2I_CONVERT;
		end case;
	end process;
	FPU_OPCODE <= fpu_opcode_s;
	
	-- INSTRUCTION TYPE DISCRIMINATOR
	discriminate_instr_type: process (opcode_s) is
	begin
		case (opcode_s) is
			when NOP =>
				op_type <= NO_TYPE;
				
			when J | JAL =>
				op_type <= J_TYPE;
				
			when ALU_I | FPU_I =>
				op_type <= R_TYPE;
				
			when LHI | LB | LH | LW | LBU | LHU | LF | LD =>
				op_type <= L_TYPE;
				
			when SB | SH | SW | SF | SD =>
				op_type <= S_TYPE;
				
			when others =>
				op_type <= I_TYPE;
		end case;
	end process;
	
	-- HAZARD CHECK PIPELINE
	hazard_pipeline: process (CLK, RST, ENB, op_type, source1_addr_s, source2_addr_s, dest_addr_s, stall_s) is
	begin
		if rising_edge(CLK) then
			if (RST = '0') then
				for i in stages_t loop
					hazard_pipe_t(i)	<= NO_TYPE;
					hazard_pipe_s1(i)	<= (others => '0');
					hazard_pipe_s2(i)	<= (others => '0');
					hazard_pipe_d(i)	<= (others => '0');
				end loop;
				
			elsif (ENB = '1') then
				if (stall_s = '1') then
					for i in DEC to DEC loop
						hazard_pipe_t(i)	<= hazard_pipe_t(i);
						hazard_pipe_s1(i)	<= hazard_pipe_s1(i);
						hazard_pipe_s2(i)	<= hazard_pipe_s2(i);
						hazard_pipe_d(i)	<= hazard_pipe_d(i);
					end loop;
					
					hazard_pipe_t(EXE)	<= NO_TYPE;
					hazard_pipe_s1(EXE)	<= (others => '0');
					hazard_pipe_s2(EXE)	<= (others => '0');
					hazard_pipe_d(EXE)	<= (others => '0');
					
					for i in MEM to WRB loop
						hazard_pipe_t(i)	<= hazard_pipe_t(i-1);
						hazard_pipe_s1(i)	<= hazard_pipe_s1(i-1);
						hazard_pipe_s2(i)	<= hazard_pipe_s2(i-1);
						hazard_pipe_d(i)	<= hazard_pipe_d(i-1);
					end loop;
					
				else
					hazard_pipe_t(DEC)	<= op_type;
					hazard_pipe_s1(DEC)	<= source1_addr_s;
					hazard_pipe_s2(DEC)	<= source2_addr_s;
					hazard_pipe_d(DEC)	<= dest_addr_s;
					for i in EXE to WRB loop
						hazard_pipe_t(i)	<= hazard_pipe_t(i-1);
						hazard_pipe_s1(i)	<= hazard_pipe_s1(i-1);
						hazard_pipe_s2(i)	<= hazard_pipe_s2(i-1);
						hazard_pipe_d(i)	<= hazard_pipe_d(i-1);
					end loop;
				end if;
			end if;
		end if;
	end process;
	
	-- FORWRDING CHECK
	-- Forwarding is checked at the earliest possible occasion (DECODE stage, if forwarding is not possible, stalling is employed).
	-- The forwarding target instruction type is checked to see whether one or more source registers are employed, then the source register(s)
	-- is/are checked against the destination register(s) of the following instructions, but only if the following instruction types
	-- require a destination register (in most cases).
	target_has_s1		<= '1' when (hazard_pipe_t(DEC) = R_TYPE or hazard_pipe_t(DEC) = I_TYPE)	else '0';
	target_has_s2		<= '1' when (hazard_pipe_t(DEC) = R_TYPE)									else '0';
	exe_source_has_d	<= '1' when not(hazard_pipe_t(EXE) = J_TYPE	or hazard_pipe_t(EXE) = S_TYPE)	else '0';
	mem_source_has_d	<= '1' when not(hazard_pipe_t(MEM) = J_TYPE	or hazard_pipe_t(MEM) = S_TYPE)	else '0';
	wrb_source_has_d	<= '1' when not(hazard_pipe_t(WRB) = J_TYPE	or hazard_pipe_t(WRB) = S_TYPE)	else '0';
	exe_can_forward_s1	<= '1' when (hazard_pipe_s1(DEC) = hazard_pipe_d(EXE))						else '0';
	mem_can_forward_s1	<= '1' when (hazard_pipe_s1(DEC) = hazard_pipe_d(MEM))						else '0';
	wrb_can_forward_s1	<= '1' when (hazard_pipe_s1(DEC) = hazard_pipe_d(WRB))						else '0';
	exe_can_forward_s2	<= '1' when (hazard_pipe_s2(DEC) = hazard_pipe_d(EXE))						else '0';
	mem_can_forward_s2	<= '1' when (hazard_pipe_s2(DEC) = hazard_pipe_d(MEM))						else '0';
	wrb_can_forward_s2	<= '1' when (hazard_pipe_s2(DEC) = hazard_pipe_d(WRB))						else '0';
	
	---- S1
	X2D_FORWARD_S1_EN	<= target_has_s1 and exe_source_has_d and exe_can_forward_s1;
	M2D_FORWARD_S1_EN	<= target_has_s1 and exe_source_has_d and mem_can_forward_s1;
	W2D_FORWARD_S1_EN	<= target_has_s1 and exe_source_has_d and wrb_can_forward_s1;
	---- S2
	X2D_FORWARD_S2_EN	<= target_has_s2 and exe_source_has_d and exe_can_forward_s2;
	M2D_FORWARD_S2_EN	<= target_has_s2 and exe_source_has_d and mem_can_forward_s2;
	W2D_FORWARD_S2_EN	<= target_has_s2 and exe_source_has_d and wrb_can_forward_s2;
	
	-- STALL CHECK
	-- Stall occurs in the particular case in which a source register requires data that has not been fetched from the main memory yet, i.e. if an instruction in the
	-- DECODE stage requires the destination of a load-type operation in the EXECUTION stage.
	-- In this case, the previous stages are disabled (with the exception of the RF in the DECODE stage) for 1 clock cycle, after which forwarding is possible.
	exe_source_is_load	<= '1' when (hazard_pipe_t(EXE) = L_TYPE) else '0';
	stall_s				<= (target_has_s1 or target_has_s2) and exe_source_is_load and (exe_can_forward_s1 or exe_can_forward_s2);
	STALL				<= stall_s;
	
end architecture;
