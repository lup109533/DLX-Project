library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.DLX_globals.all;
use work.test_instructions.all;

entity INSTR_CONVERTER is
	port (
		INSTR_IN	: in	
	);
end entity;